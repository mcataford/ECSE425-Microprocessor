library IEEE;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity CPU_tb is
end entity;

architecture CPU_tst of CPU_tb is

begin

end architecture;