library IEEE;

use ieee.std_logic_1164.all;

entity EX_STAGE is

port(

A,B,I,Ins,PC: in std_logic_vector(31 downto 0);
BRANCH: out std_logic;
R,B,Ins: out std_logic_vector(31 downto 0)

);

end entity;

architecture EX_STAGE_Impl is EX_STAGE is

begin



end architecture;