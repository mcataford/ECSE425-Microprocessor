library IEEE;

use ieee.std_logic_1164.all;

entity MEM_STAGE is

	port ();

end entity;

architecture MEM_STAGE_Impl of MEM_STAGE is

begin

end architecture;