library IEEE;

use ieee.std_logic_1164.all;

entity ALU is

end entity;

architecture ALU_impl of ALU is

begin

end architecture;