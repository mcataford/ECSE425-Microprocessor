library IEEE;

use ieee.std_logic_1164.all;

entity MICROPROCESSOR is

end entity;

architecture MICROPROCESSOR_Impl of MICROPROCESSOR is

begin

end architecture;